`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/07/11 10:10:03
// Design Name: 
// Module Name: uart_rx
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module uart_rx(
    input clk,
    input rst_n,
    input rx,
    output reg [7:0]data_out,
    output reg valid            //���ݽ������ʹ���ź�
    );
    
parameter SYSCLKHZ = 125_000_000;   //ϵͳʱ��
parameter BAUD = 115200;    //������
parameter DELAY = SYSCLKHZ/BAUD;    //����1bit����ʱ����

parameter IDLE = 4'b0001;
parameter START = 4'b0010;
parameter RESEV = 4'b0100;  //8bit���ݽ���
parameter STOP = 4'b1000;   //ֹͣλ

reg [11:0]cnt;
reg [3:0]cnt_bit;
reg [1:0]rx_temp;       //����½���
reg [3:0]state_c,state_n;

wire idl2s1_start ;
wire s12s2_start  ;
wire s22s3_start  ;
wire s32idl_start  ;

//��һ�Σ�ͬ��ʱ��alwaysģ�飬��ʽ��������̬�Ĵ���Ǩ�Ƶ���̬�Ĵ���(������ģ�
always@(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        state_c <= IDLE;
    end
    else begin
        state_c <= state_n;
    end
end

//�ڶ��Σ�����߼�alwaysģ�飬����״̬ת�������ж�
always@(*)begin
    case(state_c)
        IDLE:begin
            if(idl2s1_start)begin
                state_n = START;
            end
            else begin
                state_n = state_c;
            end
            end
        START:begin
            if(s12s2_start)begin
                state_n = RESEV;
            end
            else begin
                state_n = state_c;
            end
            end
        RESEV:begin
            if(s22s3_start)begin
                state_n = STOP;
            end
            else begin
                state_n = state_c;
            end
            end
        STOP:begin
            if(s32idl_start)begin
                state_n = IDLE;
            end
            else begin
                state_n = state_c;
            end
            end
        default:begin
            state_n = IDLE;
        end
    endcase
end

//�����Σ����ת������
assign idl2s1_start  = state_c==IDLE && rx_temp==2'b10;
assign s12s2_start = state_c==START  && cnt>=DELAY-1;
assign s22s3_start = state_c==RESEV  && cnt_bit==8 && cnt>=DELAY-1;
assign s32idl_start  = state_c==STOP && rx_temp==2'b11 || cnt>=DELAY-1;

//���ĶΣ�ͬ��ʱ��alwaysģ�飬��ʽ�������Ĵ�����������ж�������
always  @(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        cnt <=0;      //��ʼ��
        cnt_bit <=0;
        rx_temp <=0;
        data_out <=0;
        valid <=0;
    end
    else begin
        case(state_c)
            IDLE:begin
                cnt <=1'b0;
                cnt_bit <=1'b0;
                rx_temp <={rx_temp[0],rx};
                data_out <=data_out;
                valid <=1'b0;
            end
            START:begin
                if(cnt >= DELAY-1)
                    cnt <= 0;
                else
                    cnt <= cnt+1;
                cnt_bit<=0;
                data_out<=data_out;
                valid<=0;
            end
            RESEV:begin
                if(cnt>=DELAY-1)
                    cnt<=0;
                else
                    cnt<=cnt+1;
                if(cnt==(DELAY>>1))begin
                    cnt_bit<=cnt_bit+1;
                    data_out<={rx,data_out[7:1]};
                end
                else begin
                    cnt_bit <= cnt_bit;
                    data_out <= data_out;
                end
                valid<=0;
                rx_temp<={rx_temp[0],rx};
            end
            STOP:begin
                if(cnt>=DELAY-1)
                    cnt<=0;
                else
                    cnt<=cnt+1;
                rx_temp<={rx_temp[0],rx};
                data_out <= data_out;
                cnt_bit <= 0;
                if(cnt==0)
                    valid<=1;
                else
                    valid<=0;
            end
            default:begin
                cnt <=1'b0;
                cnt_bit <=1'b0;
                rx_temp <={rx_temp[0],rx};
                data_out <=data_out;
                valid <=1'b0;
            end
        endcase
    end
end
endmodule
